module frame(
	input  [64:0] frame,
	output [64:0] byte_to_seek_to
)

